LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE std.textio.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_beh IS
END tb_beh;
 
ARCHITECTURE behavior OF tb_beh IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT DCT_str
    PORT(
         Clk : IN  std_logic;
         Start : IN  std_logic;
         Din : IN  integer;
         Done : OUT  std_logic;
         Dout : OUT  integer
        );
    END COMPONENT;
    

   --Inputs
   signal Clk : std_logic := '0';
   signal Start : std_logic := '0';
   signal Din : integer := 0;

 	--Outputs
   signal Done : std_logic;
   signal Dout : integer;

   -- Clock period definitions
   constant Clk_period : time := 68 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: DCT_str PORT MAP (
          Clk => Clk,
          Start => Start,
          Din => Din,
          Done => Done,
          Dout => Dout
        );

   -- Clock process definitions
   Clk_process :process
   begin
		Clk <= '0';
		wait for Clk_period/2;
		Clk <= '1';
		wait for Clk_period/2;
   end process;


    Start <= '0' after 0 ns,
             '1' after 50 ns,
             '0' after 100 ns;


   -- Stimulus process
   stim_proc: process
   
		          variable stringbuff : LINE;
					 variable a:integer:= 1;
					 
                type RF is array ( 0 to 7, 0 to 7 ) of INTEGER;
                variable Temp   :  RF;
                variable Result :  RF;

    begin
                Temp := (
                    (49980,49980,49980,49980,49980,49980,49980,49980),
				    (-15045,-15045,-15045,-15045,-15045,-15045,-15045,-15045),
				    (87465,87465,87465,87465,87465,87465,87465,87465),
				    (-11220,-11220,-11220,-11220,-11220,-11220,-11220,-11220),
				    (51000,51000,51000,51000,51000,51000,51000,51000),
				    (34935,34935,34935,34935,34935,34935,34935,34935),
				    (20145,20145,20145,20145,20145,20145,20145,20145),
				    (37740,37740,37740,37740,37740,37740,37740,37740)
				  );
				  
				 Result := (
				      (34636140,-7147140,8946420,-649740,5747700,1549380,4048380,2848860),
                      (-10426185,    2151435,    -2693055,   195585,    -1730175,    -466395,    -1218645,    -857565),
                      (60613245,    -12507495,    15656235,  -1137045,  10058475,    2711415,    7084665,    4985505),
                      (-7775460,    1604460,    -2008380,    145860,    -1290300,    -347820,    -908820,    -639540),
                      (35343000,    -7293000,    9129000,    -663000,    5865000,    1581000,    4131000,    2907000),
                      (24209955,    -4995705,    6253365,    -454155,    4017525,    1082985,    2829735,    1991295),
                      (13960485,    -2880735,    3605955,    -261885,    2316675,    624495,    1631745,    1148265),
                      (26153820,    -5396820,    6755460,    -490620,    4340100,    1169940,    3056940,    2151180)
                  );
        
		       	WRITE (stringbuff, string'("Starts Structural Simulation at "));
		      	WRITE (stringbuff, now);
			    WRITELINE (output, stringbuff);
                ---------------------------------
                --      Handshaking/synchronizing
                ---------------------------------
                wait until Start =  '1';
                
                ---------------------------------
                --      Feed Data -- Sandwich Case
                ---------------------------------
                for i in 0 to 7 loop
                    wait until Clk = '1';
                    Din <= 255;
                end loop;
                
                for i in 0 to 4 loop
                    for j in 0 to 7 loop
                        wait until Clk = '1';
                        Din <= 0;
                    end loop;
                end loop;
                
                for i in 0 to 1 loop
                    for j in 0 to 7 loop
                        wait until Clk = '1';
                        Din <= 255;
                    end loop;
                end loop;                
                

				-- continue feeding in rest of sandwich

                ---------------------------------
                --      Handshaking/synchronizing
                ---------------------------------
                wait until Done = '1';
				wait for 5 ns;
                wait until Clk = '1' AND Clk'EVENT; 

				--------------------------------
				--      Verify
				--------------------------------
				
                for i in 0 to 7 loop
                    for j in 0 to 7 loop
                        wait until Clk = '1';
                        assert Dout = Result(i,j) report "Not Equal" SEVERITY WARNING;
                    end loop;
                end loop;
                	
				-- for each clock cycle now, start comparing values
				WRITE (stringbuff, string'("Verification completed. Simulation Ends at "));
				WRITE (stringbuff, now);
				WRITELINE (output, stringbuff);
				wait;
        end process;

END;
